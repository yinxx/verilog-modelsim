module decoder_4_12
	(
		input wire [3:0] a,
		output reg [11:0] y
	);

	// Body
	always @*
		case (a)
			4'b0000: y = 12'b000000000000;
			4'b0001: y = 12'b000000000001;
			4'b0010: y = 12'b000000000010;
			4'b0011: y = 12'b000000000100;
			4'b0100: y = 12'b000000001000;
			4'b0101: y = 12'b000000010000;
			4'b0110: y = 12'b000000100000;
			4'b0111: y = 12'b000001000000;
			4'b1000: y = 12'b000010000000;
			4'b1001: y = 12'b000100000000;
			4'b1010: y = 12'b001000000000;
			4'b1011: y = 12'b010000000000;
			4'b1100: y = 12'b100000000000;
			default: y = 12'b000000000000;
		endcase

endmodule
