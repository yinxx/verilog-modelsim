`timescale 1 ns/10 ps

module simplified_fp_greater_than_tb;
	// Signal declaration
	reg [12:0] a_test, b_test;
	wire gt_test;

	// Instantiate the circuit under test
	simplified_fp_greater_than uut
		(.a(a_test), .b(b_test), .gt(gt_test));
	
	// Test vector generator
	initial
	begin
		// Group 1
		// a = +0.68E3, b = +0.86E3 
		a_test = 13'b0101010101010;
		b_test = 13'b0101011010111;
		# 200;
		// a = -0.68E3, b = +0.86E3
		a_test = 13'b1101010101010;
		b_test = 13'b0101011010111;
		# 200;
		// a = +0.68E3, b = -0.86E3
		a_test = 13'b0101010101010;
		b_test = 13'b1101011010111;
		# 200;
		// a = -0.68E3, b = -0.86E3
		a_test = 13'b1101010101010;
		b_test = 13'b1101011010111;
		# 200;
		
		// Group 2		
		// a = +0.86E3, b = +0.68E3 
		a_test = 13'b0101011010111;
		b_test = 13'b0101010101010;
		# 200;
		// a = -0.86E3, b = +0.68E3
		a_test = 13'b1101011010111;
		b_test = 13'b0101010101010;
		# 200;
		// a = +0.86E3, b = -0.68E3
		a_test = 13'b0101011010111;
		b_test = 13'b1101010101010;
		# 200;
		// a = -0.86E3, b = -0.68E3
		a_test = 13'b1101011010111;
		b_test = 13'b1101010101010;
		# 200;
		
		// Group 3
		// a = +0.68E4, b = +0.86E3
		a_test = 13'b0110111010100;
		b_test = 13'b0101011010111;
		# 200;
		// a = -0.68E4, b = +0.86E3
		a_test = 13'b1110111010100;
		b_test = 13'b0101011010111;
		# 200;
		// a = +0.68E4, b = -0.86E3
		a_test = 13'b0110111010100;
		b_test = 13'b1101011010111;
		# 200;
		// a = -0.68E4, b = -0.86E3
		a_test = 13'b1110111010100;
		b_test = 13'b1101011010111;
		# 200;
		
		// Group 4 
		// a = +0.68E3, b = +0.86E4
		a_test = 13'b0101010101010;
		b_test = 13'b0111010000110;
		# 200;
		// a = -0.68E3, b = +0.86E4
		a_test = 13'b1101010101010;
		b_test = 13'b0111010000110;
		# 200;
		// a = +0.68E3, b = -0.86E4
		a_test = 13'b0101010101010;
		b_test = 13'b1111010000110;
		# 200;
		// a = -0.68E3, b = -0.86E4
		a_test = 13'b1101010101010;
		b_test = 13'b1111010000110;
		# 200;
		
		// Group 5
		// a = +0.68E0, b = +0.86E0
		a_test = 13'b0000010101110;
		b_test = 13'b0000011011100;
		# 200;
		// a = +0.68E0, b = -0.86E0
		a_test = 13'b0000010101110;
		b_test = 13'b1000011011100;
		# 200;

		// Group 6
		// a = +0.68E0, b = +0.68E0
		a_test = 13'b0000010101110;
		b_test = 13'b0000010101110;
		# 200;
		// a = -0.68E0, b = -0.68E0
		a_test = 13'b1000010101110;
		b_test = 13'b1000010101110;
		# 200;

		// Group 7
		// a = +0.00E0, b = +0.00E0
		a_test = 13'b0000000000000;
		b_test = 13'b0000000000000;
		# 200;
		// a = +0.00E0, b = -0.00E0
		a_test = 13'b0000000000000;
		b_test = 13'b1000000000000;
		# 200;
		
		// Stop simulation
		$stop;
	end
	
endmodule
