module fp_to_int_tb;
	// Signal declaration
	reg [12:0] fp_in_test;
	wire [7:0] int_out_test;
	wire uf_test, of_test;
	
	// Instantiate the circuit under test
	fp_to_int uut 
		(.fp_in(fp_in_test), .int_out(int_out_test), 
		.uf(uf_test), . of(of_test));
	
	// Test vector generator
	initial
	begin
		fp_in_test = 13'b0000000000000;	// +0.00000000 * 2^0 (+0)
		# 200;
		fp_in_test = 13'b1000000000000;	// -0.00000000 * 2^0 (-0)
		# 200;
		fp_in_test = 13'b0000010000000;	// +0.10000000 * 2^0 (+0.5)
		# 200;
		fp_in_test = 13'b1000010000000;	// -0.10000000 * 2^0 (-0.5)
		# 200;
		fp_in_test = 13'b0000011111111;	// +0.11111111 * 2^0 (+0.999)
		# 200;
		fp_in_test = 13'b1000011111111;	// -0.11111111 * 2^0 (-0.999)
		# 200;
		fp_in_test = 13'b0000110000000;	// +0.10000000 * 2^1 (+1)
		# 200;
		fp_in_test = 13'b1000110000000;	// -0.10000000 * 2^1 (-1)
		# 200;
		fp_in_test = 13'b0000111110000;	// +0.11110000 * 2^1 (+1.875)
		# 200;
		fp_in_test = 13'b1000111110000;	// -0.11110000 * 2^1 (-1.875)
		# 200;
		fp_in_test = 13'b0001010000000;	// +0.10000000 * 2^2 (+2)
		# 200;
		fp_in_test = 13'b1001010000000;	// -0.10000000 * 2^2 (-2)
		# 200;
		fp_in_test = 13'b0011010010000;	// +0.10010000 * 2^6 (+36)
		# 200;
		fp_in_test = 13'b1011010010000;	// -0.10010000 * 2^6 (-36)
		# 200;
		fp_in_test = 13'b0011111111110;	// +0.11111110 * 2^7 (+127)
		# 200;
		fp_in_test = 13'b1011111111110;	// -0.11111110 * 2^7 (-127)
		# 200;
		fp_in_test = 13'b0100010000000;	// +0.10000000 * 2^8 (+128)
		# 200;
		fp_in_test = 13'b1100010000000;	// -0.10000000 * 2^8 (-128)
		# 200;
		fp_in_test = 13'b0111111111111;	// +0.11111111 * 2^15 (+32460)
		# 200;
		fp_in_test = 13'b1111111111111;	// -0.11111111 * 2^15 (-32460)
		# 200;
		
		// Stop simulation
		$stop;
	end
	
endmodule
